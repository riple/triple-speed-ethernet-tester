-- Copyright (C) 1991-2011 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 10.1 Build 197 01/19/2011 Service Pack 1 SJ Full Version
-- Created on Mon Apr 25 11:17:21 2011

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY bwp_fsm IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        test_start : IN STD_LOGIC := '0';
        buffer_full : IN STD_LOGIC := '0';
        buffer_half : IN STD_LOGIC := '0';
        buffer_empty : IN STD_LOGIC := '0';
        duty_reached : IN STD_LOGIC := '0';
        cycle_reached : IN STD_LOGIC := '0';
        burst_test : IN STD_LOGIC := '0';
        burst_disabled : IN STD_LOGIC := '0';
        burst_once : IN STD_LOGIC := '0';
        buffer_ovfl : IN STD_LOGIC := '0';
        wait_once : IN STD_LOGIC := '0';
        external_int : IN STD_LOGIC := '0';
        state_ff : OUT STD_LOGIC;
        state_br : OUT STD_LOGIC;
        state_fh : OUT STD_LOGIC;
        state_sr : OUT STD_LOGIC;
        state_ti : OUT STD_LOGIC
    );
END bwp_fsm;

ARCHITECTURE BEHAVIOR OF bwp_fsm IS
    TYPE type_fstate IS (TEST_IDLE,FILL_FULL,BURST_RATE,FILL_HALF,SPACED_RATE);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
    SIGNAL reg_state_ff : STD_LOGIC := '0';
    SIGNAL reg_state_br : STD_LOGIC := '0';
    SIGNAL reg_state_fh : STD_LOGIC := '0';
    SIGNAL reg_state_sr : STD_LOGIC := '0';
    SIGNAL reg_state_ti : STD_LOGIC := '0';
BEGIN
    PROCESS (clock,reset,reg_fstate)
    BEGIN
        IF (reset='1') THEN
            fstate <= TEST_IDLE;
        ELSIF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,test_start,buffer_full,buffer_half,buffer_empty,duty_reached,cycle_reached,burst_test,burst_disabled,burst_once,buffer_ovfl,wait_once,external_int,reg_state_ff,reg_state_br,reg_state_fh,reg_state_sr,reg_state_ti)
    BEGIN
        reg_state_ff <= '0';
        reg_state_br <= '0';
        reg_state_fh <= '0';
        reg_state_sr <= '0';
        reg_state_ti <= '0';
        state_ff <= '0';
        state_br <= '0';
        state_fh <= '0';
        state_sr <= '0';
        state_ti <= '0';
        CASE fstate IS
            WHEN TEST_IDLE =>
                IF ((((test_start = '1') AND (burst_test = '1')) AND NOT((cycle_reached = '1')))) THEN
                    reg_fstate <= FILL_FULL;
                ELSIF (((test_start = '1') AND NOT((burst_test = '1')))) THEN
                    reg_fstate <= SPACED_RATE;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= TEST_IDLE;
                END IF;

                reg_state_ti <= '1';
            WHEN FILL_FULL =>
                IF ((((((buffer_full = '1') AND (buffer_ovfl = '1')) AND NOT((burst_disabled = '1'))) AND NOT((cycle_reached = '1'))) AND NOT((wait_once = '1')))) THEN
                    reg_fstate <= BURST_RATE;
                ELSIF (((((buffer_full = '1') AND (burst_disabled = '1')) AND NOT((cycle_reached = '1'))) AND NOT((wait_once = '1')))) THEN
                    reg_fstate <= SPACED_RATE;
                ELSIF (((((buffer_full = '1') AND (buffer_ovfl = '1')) AND (cycle_reached = '1')) AND NOT((wait_once = '1')))) THEN
                    reg_fstate <= TEST_IDLE;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= FILL_FULL;
                END IF;

                reg_state_ff <= '1';
            WHEN BURST_RATE =>
                IF ((((buffer_empty = '1') AND NOT((burst_once = '1'))) AND NOT((burst_disabled = '1')))) THEN
                    reg_fstate <= FILL_HALF;
                ELSIF (((burst_disabled = '1') OR ((buffer_empty = '1') AND (burst_once = '1')))) THEN
                    reg_fstate <= SPACED_RATE;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= BURST_RATE;
                END IF;

                reg_state_br <= '1';
            WHEN FILL_HALF =>
                IF ((buffer_half = '1')) THEN
                    reg_fstate <= SPACED_RATE;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= FILL_HALF;
                END IF;

                reg_state_fh <= '1';
            WHEN SPACED_RATE =>
                IF ((((((duty_reached = '1') AND (burst_test = '1')) AND NOT((burst_disabled = '1'))) AND NOT((burst_once = '1'))) OR (((external_int = '1') AND (burst_test = '1')) AND (burst_once = '1')))) THEN
                    reg_fstate <= FILL_FULL;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= SPACED_RATE;
                END IF;

                reg_state_sr <= '1';
            WHEN OTHERS => 
                reg_state_ff <= 'X';
                reg_state_br <= 'X';
                reg_state_fh <= 'X';
                reg_state_sr <= 'X';
                reg_state_ti <= 'X';
                report "Reach undefined state";
        END CASE;
        state_ff <= reg_state_ff;
        state_br <= reg_state_br;
        state_fh <= reg_state_fh;
        state_sr <= reg_state_sr;
        state_ti <= reg_state_ti;
    END PROCESS;
END BEHAVIOR;
